set_property PACKAGE_PIN W5 [get_ports clock]							
	set_property IOSTANDARD LVCMOS33 [get_ports clock]
	create_clock -add -name sys_clk_pin -period 10.00 -waveform {0 5} [get_ports clock]
	
set_property PACKAGE_PIN U18 [get_ports clear]						
    set_property IOSTANDARD LVCMOS33 [get_ports clear]
    
set_property PACKAGE_PIN V17 [get_ports stop]					
        set_property IOSTANDARD LVCMOS33 [get_ports stop]
    
set_property PACKAGE_PIN W7 [get_ports {a_to_g[0]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {a_to_g[0]}]
set_property PACKAGE_PIN W6 [get_ports {a_to_g[1]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {a_to_g[1]}]
set_property PACKAGE_PIN U8 [get_ports {a_to_g[2]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {a_to_g[2]}]
set_property PACKAGE_PIN V8 [get_ports {a_to_g[3]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {a_to_g[3]}]
set_property PACKAGE_PIN U5 [get_ports {a_to_g[4]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {a_to_g[4]}]
set_property PACKAGE_PIN V5 [get_ports {a_to_g[5]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {a_to_g[5]}]
set_property PACKAGE_PIN U7 [get_ports {a_to_g[6]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {a_to_g[6]}]

set_property PACKAGE_PIN U2 [get_ports {an[0]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {an[0]}]
set_property PACKAGE_PIN U4 [get_ports {an[1]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {an[1]}]
set_property PACKAGE_PIN V4 [get_ports {an[2]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {an[2]}]
set_property PACKAGE_PIN W4 [get_ports {an[3]}]					
	set_property IOSTANDARD LVCMOS33 [get_ports {an[3]}]